module vram_ctrl(
						input wire clk, reset,
						
						//From video sync
						input wire [9:0] pixel_x, pixel_y,
						input wire p_tick,
						
						//Memory interface to VGA read
						output wire [7:0] vga_rd_data,
						
						//Memory interface to GPU
						input wire cpu_mem_wr, cpu_mem_rd,
						input wire [18:0] cpu_addr,
						input wire [7:0] cpu_wr_data,
						output wire [7:0] cpu_rd_data,
						
						//To and From SRAM
						output wire [17:0] sram_addr,
						inout [15:0] sram_dq,
						output sram_ce_n, sram_oe_n, sram_wr_n,
						output sram_lb_n, sram_ub_n
						);
						
//States
localparam [2:0] idle = 3'd0,
					  waitr = 3'd1,
					  rd = 3'd2,
					  fetch = 3'd3,
					  waitw = 3'd4,
					  wr = 3'd5;
					  
//Signal declarations
reg [2:0] state_reg, state_next;
reg [7:0] vga_rd_data_reg;
reg [18:0] cpu_addr_reg, cpu_addr_next;
wire [18:0] mem_addr;
wire [18:0] y_offset, vga_addr; //why offset?
reg [7:0] cpu_rd_data_reg, cpu_rd_data_next;
reg [7:0] wr_data_reg, wr_data_next;
reg we_n_reg;
wire we_n_next;
wire [7:0] byte_from_sram;
wire vga_cycle;

//what is p-tick doing?
//p-tick is asserted every 2 clock cycles

//*****************************************************
// VGA port SRAM read operation
//*****************************************************

//VGA Port reads SRAM contunuously

always@(posedge clk) begin
	
	if (vga_cycle)	vga_rd_data_reg <= byte_from_sram;
		
end

assign y_offset = {1'd0, pixel_y[8:0], 9'd0} + {3'd0, pixel_y[8:0], 7'd0};
assign vga_addr = y_offset + pixel_x;
assign vga_rd_data = vga_rd_data_reg;

//*****************************************************
// CPU port SRAM read-write operation
//*****************************************************

assign cpu_rd_data= cpu_rd_data_reg; 
// FSMD state & data registers
always @(posedge clk, posedge reset) begin 
	if (reset) begin
		state_reg <= idle;
		cpu_addr_reg <= 0;
		wr_data_reg <= 0;
		cpu_rd_data_reg <= 0;
	end
	else begin
		state_reg <= state_next;
		cpu_addr_reg <= cpu_addr_next;
		wr_data_reg <= wr_data_next;
		cpu_rd_data_reg <= cpu_rd_data_next; we_n_reg <= we_n_next;
	end
end
// FSMD next-state logic	
always@(*) begin
	state_next = state_reg;
	cpu_addr_next = cpu_addr_reg;
	wr_data_next = wr_data_reg;
	cpu_rd_data_next = cpu_rd_data_reg;

	case (state_reg)
		idle:
			if (cpu_mem_wr)
			begin
				
					cpu_addr_next = cpu_addr;
					cpu_addr_next = wr_data_next;
					
					if (vga_cycle) 
						state_next = wr;
					else 
						state_next = waitw;
			end	
			else if (cpu_mem_rd) begin
			
					if (vga_cycle)
						state_next = rd;
					else begin
						state_next = waitr;
						cpu_rd_data_next = byte_from_sram;
					end
				end
	
		rd: begin
				cpu_rd_data_next = byte_from_sram; 
				state_next = fetch;
			end
		waitr:
			state_next = fetch;
		
		fetch:
			state_next = idle;
		
		waitw:
			state_next = wr;
		
		wr: 
			state_next = idle;
			
	endcase
end


// look-ahead output
assign we_n_next = (state_next==wr) ? 1'b0: 1'b1;


//*****************************************************
// SRAM interface signals
//*****************************************************

// configure SRAM as 512K-by-8
assign mem_addr = vga_cycle ? vga_addr:
													((~we_n_reg) ? cpu_addr_reg:cpu_addr);

assign sram_addr = mem_addr [18:1];
assign sram_lb_n = (~mem_addr [0]) ? 1'b0: 1'b1;
assign sram_ub_n = (mem_addr [0]) ? 1'b0: 1'b1;
assign sram_ce_n = 1'b0;
assign sram_oe_n = 1'b0;
assign sram_we_n = we_n_reg;
assign sram_dq = (~we_n_reg)? {wr_data_reg, wr_data_reg}: 16'bz;

// LSB control lb ub
assign byte_from_sram = mem_addr [0] ? sram_dq [15:8]: sram_dq [7:0];

endmodule			
			
			

